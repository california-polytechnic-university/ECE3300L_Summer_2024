`timescale 1ns / 1ps

module tb_Decoder4x16;

reg [3:0] SW;  // 4 input switches
wire [15:0] LED;  // 16 output LEDs

// Instantiate the Decoder4x16 module
Decoder4x16 uut (
    .SW(SW),
    .LED(LED)
);

initial begin
    // Apply test vectors
    SW = 4'b0000; #10;
    SW = 4'b0001; #10;
    SW = 4'b0010; #10;
    SW = 4'b0011; #10;
    SW = 4'b0100; #10;
    SW = 4'b0101; #10;
    SW = 4'b0110; #10;
    SW = 4'b0111; #10;
    SW = 4'b1000; #10;
    SW = 4'b1001; #10;
    SW = 4'b1010; #10;
    SW = 4'b1011; #10;
    SW = 4'b1100; #10;
    SW = 4'b1101; #10;
    SW = 4'b1110; #10;
    SW = 4'b1111; #10;
    
    // End simulation
    $stop;
end

endmodule
