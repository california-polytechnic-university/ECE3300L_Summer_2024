`timescale 1ns / 1ps
module decoder_4x16(
     input [3:0] sw,
     output reg [15:0] led

    );
    always @(*) begin
        case (sw)
            4'b0000: led = 16'b0000000000000001;
            4'b0001: led = 16'b0000000000000010;
            4'b0010: led = 16'b0000000000000100;
            4'b0011: led = 16'b0000000000001000;
            4'b0100: led = 16'b0000000000010000;
            4'b0101: led = 16'b0000000000100000;
            4'b0110: led = 16'b0000000001000000;
            4'b0111: led = 16'b0000000010000000;
            4'b1000: led = 16'b0000000100000000;
            4'b1001: led = 16'b0000001000000000;
            4'b1010: led = 16'b0000010000000000;
            4'b1011: led = 16'b0000100000000000;
            4'b1100: led = 16'b0001000000000000;
            4'b1101: led = 16'b0010000000000000;
            4'b1110: led = 16'b0100000000000000;
            4'b1111: led = 16'b1000000000000000;
            default: led = 16'b0000000000000000;
        endcase
    end
    
endmodule
