`timescale 1ns / 1ps

module mux4x1_tb;
    
    reg [13:0] sw;
    wire [2:0] led;
    
    topmod dut (
        .top_sw(sw),
        .top_led(led)
    );
    
    
initial 
   begin
        //start position for test
            sw = 14'b0000_0000_0000_00;
            
            //sel = 00
            #10
            sw = 14'b0000_0000_0000_00;
            #10
            sw = 14'b0000_0000_0001_00;
            #10
            sw = 14'b0000_0001_0000_00;
            #10
            sw = 14'b0001_0000_0000_00;
            #10
            sw = 14'b0001_0001_0000_00;
            #10
            sw = 14'b0000_0001_0001_00;
            #10
            sw = 14'b0001_0000_0001_00;
            #10
            sw = 14'b0001_0001_0001_00;
            
            //sel 01
            #10
            sw = 14'b0000_0000_0000_01;
            #10
            sw = 14'b0000_0000_0010_01;
            #10
            sw = 14'b0000_0010_0000_01;
            #10
            sw = 14'b0010_0000_0000_01;
            #10
            sw = 14'b0010_0010_0000_01;
            #10
            sw = 14'b0000_0010_0010_01;
            #10
            sw = 14'b0010_0000_0010_01;
            #10
            sw = 14'b0010_0010_0010_01;
            
            //sel 10
            #10
            sw = 14'b0000_0000_0000_10;
            #10
            sw = 14'b0000_0000_0100_10;
            #10
            sw = 14'b0000_0100_0000_10;
            #10
            sw = 14'b0100_0000_0000_10;
            #10
            sw = 14'b0100_0100_0000_10;
            #10
            sw = 14'b0000_0100_0100_10;
            #10
            sw = 14'b0100_0000_0100_10;
            #10
            sw = 14'b0100_0100_0100_10;
            
            //sel 11
            #10
            sw = 14'b0000_0000_0000_11;
            #10
            sw = 14'b0000_0000_1000_11;
            #10
            sw = 14'b0000_1000_0000_11;
            #10
            sw = 14'b1000_0000_0000_11;
            #10
            sw = 14'b1000_1000_0000_11;
            #10
            sw = 14'b0000_1000_1000_11;
            #10
            sw = 14'b1000_0000_1000_11;
            #10
            sw = 14'b1000_1000_1000_11;
            #10
    $finish;
   end
endmodule
