`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/11/2024 09:27:55 PM
// Design Name: 
// Module Name: testbench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module testbench();

    reg [15:0] SW;
    wire [15:0] LED;
    
switch dut(
    .SW(SW),
    .LED(LED)
);

initial begin
    SW = 16'b0000000000000000; #10;
    SW = 16'b0000000000000001; #10;
    SW = 16'b0000000000000010; #10;
    SW = 16'b0000000000000100; #10;
    SW = 16'b0000000000001000; #10;
    SW = 16'b0000000000010000; #10;
    SW = 16'b0000000000100000; #10;
    SW = 16'b0000000001000000; #10;
    SW = 16'b0000000010000000; #10;
    SW = 16'b0000000100000000; #10;
    SW = 16'b0000001000000000; #10;
    SW = 16'b0000010000000000; #10;
    SW = 16'b0000100000000000; #10;
    SW = 16'b0001000000000000; #10;
    SW = 16'b0010000000000000; #10;
    SW = 16'b0100000000000000; #10;
    SW = 16'b1000000000000000; #10;
    SW = 16'b1111111111111111; #10;
    $finish;
    end
endmodule
